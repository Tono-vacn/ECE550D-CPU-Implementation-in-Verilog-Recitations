module alu_b(data_operandA, data_operandB, ctrl_ALUopcode, ctrl_shiftamt, data_result, isNotEqual, isLessThan, overflow);
   input [31:0] data_operandA, data_operandB;
   input [4:0] ctrl_ALUopcode, ctrl_shiftamt;

   output reg [31:0] data_result;
   output reg isNotEqual, isLessThan, overflow;
	
	localparam
		AD = 5'b00000,
		SU = 5'b00001,
		AN = 5'b00010,
		OR = 5'b00011,
		SL = 5'b00100,
		SR = 5'b00101;
	
	always@(data_operandA or data_operandB or ctrl_ALUopcode or ctrl_shiftamt) begin
		case(ctrl_ALUopcode)
			AD:
				begin
					data_result = data_operandA + data_operandB;
					overflow = (data_operandA[31]&data_operandB[31]&!data_result[31])|(!data_operandA[31]&!data_operandB[31]&data_result[31]);
				end
			SU:
				begin
					data_result = data_operandA - data_operandB;
					overflow = (data_operandA[31]&!data_operandB[31]&!data_result[31])|(!data_operandA[31]&data_operandB[31]&data_result[31]);					
				end
			AN:
				begin
					data_result = data_operandA & data_operandB;
				end
			OR:
				begin
					data_result = data_operandA | data_operandB;
				end
			SL:
				begin
					data_result = data_operandA << ctrl_shiftamt;
				end
			SR:
				begin
					data_result = $signed(data_operandA) >>> ctrl_shiftamt;
				end
			default:
				begin
				end
		endcase
		
		isNotEqual <= (data_operandA != data_operandB) ? 1'b1:1'b0;
		isLessThan <= (data_operandA[31] & !data_operandB[31])|((data_operandA[31] ~^ data_operandB[31]) & data_result[31]);
			
	end
	
endmodule
