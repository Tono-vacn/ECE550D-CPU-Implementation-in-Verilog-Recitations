module rca_8(a,b,cin,sum,cout);
	input [7:0]a,b;
	input cin;
	output [7:0]sum;
	output cout;
	
	wire [6:0]out;
	
	full_adder fa0(.a(a[0]),.b(b[0]),.cin(cin),.sum(sum[0]),.cout(out[0]));
	
	generate
		genvar i;
		for(i=1;i<7;i=i+1) begin:loop_rca8
			full_adder fa(.a(a[i]),.b(b[i]),.cin(out[i-1]),.sum(sum[i]),.cout(out[i]));
		end
	endgenerate
		
	full_adder fa1(.a(a[7]),.b(b[7]),.cin(out[6]),.sum(sum[7]),.cout(cout));
endmodule



module rca_8_overflow(a,b,cin,sum,cout,of);
	input [7:0]a,b;
	input cin;
	output [7:0]sum;
	output cout;
	output of;
	
	wire [6:0]out;
	
	full_adder fa0(.a(a[0]),.b(b[0]),.cin(cin),.sum(sum[0]),.cout(out[0]));
	
	generate
		genvar i;
		for(i=1;i<7;i=i+1) begin:loop_rca8
			full_adder fa(.a(a[i]),.b(b[i]),.cin(out[i-1]),.sum(sum[i]),.cout(out[i]));
		end
	endgenerate
		
	full_adder fa1(.a(a[7]),.b(b[7]),.cin(out[6]),.sum(sum[7]),.cout(cout));
	
	xor testof(of,cout,out[6]);
endmodule